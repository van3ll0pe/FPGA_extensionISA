module CRC32();

endmodule;